import Arbitration :: *;
import ClientServer :: *;
import Cntrs :: *;
import Connectable :: *;
import FIFOF :: *;
import GetPut :: *;
import PAClib :: *;
import Vector :: *;

import Controller :: *;
import DataTypes :: *;
import DupReadAtomicCache :: *;
import InputPktHandle :: *;
import Headers :: *;
import MetaData :: *;
import PayloadConAndGen :: *;
import PrimUtils :: *;
import RetryHandleSQ :: *;
import ReqGenSQ :: *;
import ReqHandleRQ :: *;
import RespHandleSQ :: *;
import Settings :: *;
import SpecialFIFOF :: *;
import WorkCompGen :: *;
import Utils :: *;

typedef Vector#(portSz, PermCheckSrv) PermCheckSrvArbiter#(numeric type portSz);

module mkPermCheckSrvArbiter#(PermCheckSrv permCheckSrv)(PermCheckSrvArbiter#(portSz)) provisos(
    Add#(1, anysize, portSz),
    Add#(TLog#(portSz), 1, TLog#(TAdd#(portSz, 1))) // portSz must be power of 2
);
    function Bool isPermCheckReqFinished(PermCheckReq req) = True;
    function Bool isPermCheckRespFinished(Bool resp) = True;

    PermCheckSrvArbiter#(portSz) arbiter <- mkServerArbiter(
        permCheckSrv,
        isPermCheckReqFinished,
        isPermCheckRespFinished
    );
    return arbiter;
endmodule

interface DmaArbiterInsideQP;
    interface DmaReadSrv  dmaReadSrv4RQ;
    interface DmaWriteSrv dmaWriteSrv4RQ;
    interface DmaReadSrv  dmaReadSrv4SQ;
    interface DmaWriteSrv dmaWriteSrv4SQ;
endinterface

module mkDmaArbiterInsideQP#(
    DmaReadSrv  dmaReadSrv,
    DmaWriteSrv dmaWriteSrv
)(DmaArbiterInsideQP);
    FIFOF#(DmaReadReq)     dmaReadReqQ4RQ <- mkFIFOF;
    FIFOF#(DmaReadResp)   dmaReadRespQ4RQ <- mkFIFOF;
    FIFOF#(DmaWriteReq)   dmaWriteReqQ4RQ <- mkFIFOF;
    FIFOF#(DmaWriteResp) dmaWriteRespQ4RQ <- mkFIFOF;

    FIFOF#(DmaReadReq)     dmaReadReqQ4SQ <- mkFIFOF;
    FIFOF#(DmaReadResp)   dmaReadRespQ4SQ <- mkFIFOF;
    FIFOF#(DmaWriteReq)   dmaWriteReqQ4SQ <- mkFIFOF;
    FIFOF#(DmaWriteResp) dmaWriteRespQ4SQ <- mkFIFOF;

    // RQ has higher priority than SQ when issueing DMA requests
    // and receiving DMA responses.
    rule issueDmaReadReq;
        if (dmaReadReqQ4RQ.notEmpty) begin
            let rqDmaReadReq = dmaReadReqQ4RQ.first;
            dmaReadReqQ4RQ.deq;
            dmaReadSrv.request.put(rqDmaReadReq);
        end
        else if (dmaReadReqQ4SQ.notEmpty) begin
            let sqDmaReadReq = dmaReadReqQ4SQ.first;
            dmaReadReqQ4SQ.deq;
            dmaReadSrv.request.put(sqDmaReadReq);
        end
    endrule

    rule issueDmaWriteReq;
        if (dmaWriteReqQ4RQ.notEmpty) begin
            let rqDmaWriteReq = dmaWriteReqQ4RQ.first;
            dmaWriteReqQ4RQ.deq;
            dmaWriteSrv.request.put(rqDmaWriteReq);
        end
        else if (dmaWriteReqQ4SQ.notEmpty) begin
            let sqDmaWriteReq = dmaWriteReqQ4SQ.first;
            dmaWriteReqQ4SQ.deq;
            dmaWriteSrv.request.put(sqDmaWriteReq);
        end
    endrule

    rule recvDmaReadResp;
        let dmaReadResp <- dmaReadSrv.response.get;
        case (dmaReadResp.initiator)
            DMA_INIT_RQ_RD    ,
            DMA_INIT_RQ_WR    ,
            DMA_INIT_RQ_DUP_RD,
            DMA_INIT_RQ_ATOMIC: dmaReadRespQ4RQ.enq(dmaReadResp);
            default           : dmaReadRespQ4SQ.enq(dmaReadResp);
        endcase
    endrule

    rule recvDmaWriteResp;
        let dmaWriteResp <- dmaWriteSrv.response.get;
        case (dmaWriteResp.initiator)
            DMA_INIT_RQ_RD    ,
            DMA_INIT_RQ_WR    ,
            DMA_INIT_RQ_DUP_RD,
            DMA_INIT_RQ_ATOMIC: dmaWriteRespQ4RQ.enq(dmaWriteResp);
            default           : dmaWriteRespQ4SQ.enq(dmaWriteResp);
        endcase
    endrule

    interface dmaReadSrv4RQ  = toGPServer(dmaReadReqQ4RQ,  dmaReadRespQ4RQ);
    interface dmaWriteSrv4RQ = toGPServer(dmaWriteReqQ4RQ, dmaWriteRespQ4RQ);
    interface dmaReadSrv4SQ  = toGPServer(dmaReadReqQ4SQ,  dmaReadRespQ4SQ);
    interface dmaWriteSrv4SQ = toGPServer(dmaWriteReqQ4SQ, dmaWriteRespQ4SQ);
endmodule

typedef Vector#(portSz, DmaReadSrv) DmaReadSrvArbiter#(numeric type portSz);
typedef Vector#(portSz, DmaWriteSrv) DmaWriteSrvArbiter#(numeric type portSz);

module mkDmaReadSrvArbiter#(DmaReadSrv dmaReadSrv)(DmaReadSrvArbiter#(portSz)) provisos(
    Add#(1, anysize, portSz),
    Add#(TLog#(portSz), 1, TLog#(TAdd#(portSz, 1))) // portSz must be power of 2
);
    function Bool isDmaReadReqLastFrag(DmaReadReq req) = True;
    function Bool isDmaReadRespLastFrag(DmaReadResp resp) = resp.dataStream.isLast;

    DmaReadSrvArbiter#(portSz) arbiter <- mkServerArbiter(
        dmaReadSrv,
        isDmaReadReqLastFrag,
        isDmaReadRespLastFrag
    );
    return arbiter;
endmodule

module mkDmaWriteSrvArbiter#(DmaWriteSrv dmaWriteSrv)(
    DmaWriteSrvArbiter#(portSz)
) provisos(
    Add#(1, anysize, portSz),
    Add#(TLog#(portSz), 1, TLog#(TAdd#(portSz, 1))) // portSz must be power of 2
);
    function Bool isDmaWriteReqLastFrag(DmaWriteReq req) = req.dataStream.isLast;
    function Bool isDmaWriteRespLastFrag(DmaWriteResp resp) = True;

    DmaWriteSrvArbiter#(portSz) arbiter <- mkServerArbiter(
        dmaWriteSrv,
        isDmaWriteReqLastFrag,
        isDmaWriteRespLastFrag
    );
    return arbiter;
endmodule

module mkNewPendingWorkReqPipeOut#(
    PipeOut#(WorkReq) workReqPipeIn
)(PipeOut#(PendingWorkReq));
    FIFOF#(PendingWorkReq) newPendingWorkReqOutQ <- mkFIFOF;

    rule genPendingWR;
        let wr = workReqPipeIn.first;
        workReqPipeIn.deq;

        let newPendingWR = genNewPendingWorkReq(wr);
        newPendingWorkReqOutQ.enq(newPendingWR);
    endrule

    return convertFifo2PipeOut(newPendingWorkReqOutQ);
endmodule

interface SQ;
    interface DataStreamPipeOut rdmaReqDataStreamPipeOut;
    interface PipeOut#(WorkComp) workCompPipeOutSQ;
endinterface

module mkSQ#(
    Controller cntrl,
    DmaReadSrv dmaReadSrv,
    DmaWriteSrv dmaWriteSrv,
    PermCheckSrv permCheckSrv,
    PipeOut#(WorkReq) workReqPipeIn,
    RdmaPktMetaDataAndPayloadPipeOut respPktPipeOut,
    PipeOut#(WorkCompStatus) workCompStatusPipeInFromRQ
)(SQ);
    PendingWorkReqBuf pendingWorkReqBuf <- mkScanFIFOF;

    let retryHandler <- mkRetryHandleSQ(
        cntrl, pendingWorkReqBuf.fifof.notEmpty, pendingWorkReqBuf.scanCntrl
    );

    let newPendingWorkReqPiptOut <- mkNewPendingWorkReqPipeOut(workReqPipeIn);
    // let newPendingWorkReqPiptOut = genNewPendingWorkReqPipeOut(workReqPipeIn);
    let pendingWorkReqPipeOut <- mkPipeOutMux(
        pendingWorkReqBuf.scanCntrl.hasScanOut,
        pendingWorkReqBuf.scanPipeOut,
        newPendingWorkReqPiptOut
    );

    let reqGenSQ <- mkReqGenSQ(
        cntrl, dmaReadSrv, pendingWorkReqPipeOut, pendingWorkReqBuf.fifof.notEmpty
    );
    let pendingWorkReq2Q <- mkConnectPendingWorkReqPipeOut2PendingWorkReqQ(
        reqGenSQ.pendingWorkReqPipeOut, pendingWorkReqBuf.fifof
    );

    let respHandleSQ <- mkRespHandleSQ(
        cntrl,
        retryHandler,
        permCheckSrv,
        convertFifo2PipeOut(pendingWorkReqBuf.fifof),
        respPktPipeOut.pktMetaData
    );

    let payloadConsumer <- mkPayloadConsumer(
        cntrl,
        respPktPipeOut.payload,
        dmaWriteSrv,
        respHandleSQ.payloadConReqPipeOut
    );

    let workCompPipeOut <- mkWorkCompGenSQ(
        cntrl,
        payloadConsumer.respPipeOut,
        reqGenSQ.workCompGenReqPipeOut,
        respHandleSQ.workCompGenReqPipeOut,
        workCompStatusPipeInFromRQ
    );

    interface rdmaReqDataStreamPipeOut = reqGenSQ.rdmaReqDataStreamPipeOut;
    interface workCompPipeOutSQ = workCompPipeOut;
endmodule

interface RQ;
    interface DataStreamPipeOut rdmaRespDataStreamPipeOut;
    interface PipeOut#(WorkComp) workCompPipeOutRQ;
    interface PipeOut#(WorkCompStatus) workCompStatusPipeOutRQ;
endinterface

module mkRQ#(
    Controller cntrl,
    DmaReadSrv dmaReadSrv,
    DmaWriteSrv dmaWriteSrv,
    PermCheckSrv permCheckSrv,
    RecvReqBuf recvReqBuf,
    RdmaPktMetaDataAndPayloadPipeOut reqPktPipeIn
)(RQ);
    let dupReadAtomicCache <- mkDupReadAtomicCache(cntrl.cntrlStatus.getPMTU);

    let reqHandlerRQ <- mkReqHandleRQ(
        cntrl,
        dmaReadSrv,
        permCheckSrv,
        dupReadAtomicCache,
        recvReqBuf,
        reqPktPipeIn.pktMetaData
    );

    let payloadConsumer <- mkPayloadConsumer(
        cntrl,
        reqPktPipeIn.payload,
        dmaWriteSrv,
        reqHandlerRQ.payloadConReqPipeOut
    );

    let workCompGenRQ <- mkWorkCompGenRQ(
        cntrl,
        payloadConsumer.respPipeOut,
        reqHandlerRQ.workCompGenReqPipeOut
    );

    interface rdmaRespDataStreamPipeOut = reqHandlerRQ.rdmaRespDataStreamPipeOut;
    interface workCompPipeOutRQ = workCompGenRQ.workCompPipeOut;
    interface workCompStatusPipeOutRQ = workCompGenRQ.workCompStatusPipeOutRQ;
endmodule

interface QP;
    interface DataStreamPipeOut rdmaReqRespPipeOut;
    interface PipeOut#(WorkComp) workCompPipeOutRQ;
    interface PipeOut#(WorkComp) workCompPipeOutSQ;
endinterface

module mkQP#(
    Controller cntrl,
    PipeOut#(RecvReq) recvReqPipeIn,
    PipeOut#(WorkReq) workReqPipeIn,
    DmaReadSrv dmaReadSrv,
    DmaWriteSrv dmaWriteSrv,
    PermCheckSrv permCheck4RQ,
    PermCheckSrv permCheck4SQ,
    RdmaPktMetaDataAndPayloadPipeOut reqPktPipeIn,
    RdmaPktMetaDataAndPayloadPipeOut respPktPipeIn
)(QP);
    // TODO: change WR and RR queues to mkSizedFIFOF
    FIFOF#(RecvReq) recvReqQ <- mkFIFOF;
    FIFOF#(WorkReq) workReqQ <- mkFIFOF;
    mkConnection(toPut(recvReqQ), toGet(recvReqPipeIn));
    mkConnection(toPut(workReqQ), toGet(workReqPipeIn));
    let recvReqBufPipeOut = convertFifo2PipeOut(recvReqQ);
    let workReqBufPipeOut = convertFifo2PipeOut(workReqQ);
    // let recvReqBufPipeOut <- mkPipeOutBuffer(recvReqPipeIn);
    // let workReqBufPipeOut <- mkPipeOutBuffer(workReqPipeIn);

    let dmaArbiter <- mkDmaArbiterInsideQP(
        dmaReadSrv, dmaWriteSrv
    );

    let rq <- mkRQ(
        cntrl,
        dmaArbiter.dmaReadSrv4RQ,
        dmaArbiter.dmaWriteSrv4RQ,
        permCheck4RQ,
        recvReqBufPipeOut,
        reqPktPipeIn
    );

    let sq <- mkSQ(
        cntrl,
        dmaArbiter.dmaReadSrv4SQ,
        dmaArbiter.dmaWriteSrv4SQ,
        permCheck4SQ,
        workReqBufPipeOut,
        respPktPipeIn,
        rq.workCompStatusPipeOutRQ
    );
    let reqRespPipeOut <- mkFixedBinaryPipeOutArbiter(
        rq.rdmaRespDataStreamPipeOut, sq.rdmaReqDataStreamPipeOut
    );
    rule errFlush if (cntrl.cntrlStatus.isERR);
        // TODO: if pending WR queue is empty, then error flush is done
        if (!workReqQ.notEmpty && !recvReqQ.notEmpty) begin
            // Notify controller when flush done
            cntrl.errFlushDone;
            $display(
                "time=%0t:", $time,
                " error flush done, workReqQ.notEmpty=", fshow(workReqQ.notEmpty),
                ", recvReqQ.notEmpty=", fshow(recvReqQ.notEmpty)
            );
        end
    endrule

    interface rdmaReqRespPipeOut = reqRespPipeOut;
    interface workCompPipeOutRQ = rq.workCompPipeOutRQ;
    interface workCompPipeOutSQ = sq.workCompPipeOutSQ;
endmodule

typedef union tagged {
    WorkReq WR;
    RecvReq RR;
} WorkReqOrRecvReq deriving(Bits);

// TODO: check QP state when dispatching WR and RR
module mkWorkReqAndRecvReqDispatcher#(
    PipeOut#(WorkReqOrRecvReq) workReqOrRecvReqPipeIn
)(Tuple2#(Vector#(MAX_QP, PipeOut#(WorkReq)), Vector#(MAX_QP, PipeOut#(RecvReq))));
    Vector#(MAX_QP, FIFOF#(WorkReq)) workReqOutVec <- replicateM(mkFIFOF);
    Vector#(MAX_QP, FIFOF#(RecvReq)) recvReqOutVec <- replicateM(mkFIFOF);

    rule dispatchWorkReqOrRecvReq;
        case (workReqOrRecvReqPipeIn.first) matches
            tagged WR .wr: begin
                let qpIndex = getIndexQP(wr.sqpn);
                workReqOutVec[qpIndex].enq(wr);
            end
            tagged RR .rr: begin
                let qpIndex = getIndexQP(rr.sqpn);
                recvReqOutVec[qpIndex].enq(rr);
            end
        endcase
        workReqOrRecvReqPipeIn.deq;
    endrule

    return tuple2(
        map(convertFifo2PipeOut, workReqOutVec),
        map(convertFifo2PipeOut, recvReqOutVec)
    );
endmodule

interface TransportLayerRDMA;
    interface Put#(DataStream) rdmaDataStreamInput;
    interface DataStreamPipeOut rdmaDataStreamPipeOut;
    interface Server#(WorkReqOrRecvReq, WorkComp) srvWorkReqRecvReqWorkComp;
    interface MetaDataSrv srvMetaData;
endinterface

(* synthesize *)
module mkTransportLayerRDMA(TransportLayerRDMA);
    FIFOF#(DataStream) inputDataStreamQ <- mkFIFOF;
    let rdmaReqRespPipeIn = convertFifo2PipeOut(inputDataStreamQ);

    FIFOF#(WorkReqOrRecvReq) inputWorkReqOrRecvReqQ <- mkFIFOF;

    let pdMetaData  <- mkMetaDataPDs;
    let permCheckSrv <- mkPermCheckSrv(pdMetaData);
    let qpMetaData  <- mkMetaDataQPs;
    let metaDataSrv <- mkMetaDataSrv(pdMetaData, qpMetaData);

    // let qpInitAttr = QpInitAttr {
    //     qpType  : IBV_QPT_RC,
    //     sqSigAll: False
    // };
    // let qpAttrPipeOut <- mkQpAttrPipeOut;
    // let initMetaData <- mkInitMetaData(metaDataSrv, qpInitAttr, qpAttrPipeOut);

    let { workReqPipeOutVec, recvPipeOutVec } <- mkWorkReqAndRecvReqDispatcher(
        convertFifo2PipeOut(inputWorkReqOrRecvReqQ)
    );

    PermCheckSrvArbiter#(TMul#(2, MAX_QP)) permCheckSrvArbiter <- mkPermCheckSrvArbiter(permCheckSrv);

    let headerAndMetaDataAndPayloadPipeOut <- mkExtractHeaderFromRdmaPktPipeOut(
        rdmaReqRespPipeIn
    );
    let pktMetaDataAndPayloadPipeOutVec <- mkInputRdmaPktBufAndHeaderValidation(
        headerAndMetaDataAndPayloadPipeOut, qpMetaData
    );

    let dmaReadSrv  <- mkDmaReadSrv;
    let dmaWriteSrv <- mkDmaWriteSrv;
    DmaReadSrvArbiter#(MAX_QP)   dmaReadSrvVec <- mkDmaReadSrvArbiter(dmaReadSrv);
    DmaWriteSrvArbiter#(MAX_QP) dmaWriteSrvVec <- mkDmaWriteSrvArbiter(dmaWriteSrv);

    Vector#(MAX_QP, DataStreamPipeOut)    qpDataStreamPipeOutVec = newVector;
    Vector#(MAX_QP, PipeOut#(WorkComp)) qpRecvWorkCompPipeOutVec = newVector;
    Vector#(MAX_QP, PipeOut#(WorkComp)) qpSendWorkCompPipeOutVec = newVector;

    for (Integer idx = 0; idx < valueOf(MAX_QP); idx = idx + 1) begin
        let permCheck4RQ = permCheckSrvArbiter[2 * idx];
        let permCheck4SQ = permCheckSrvArbiter[2 * idx + 1];

        IndexQP qpIndex = fromInteger(idx);
        let cntrl = qpMetaData.getCntrlByIndexQP(qpIndex);
        let qp <- mkQP(
            cntrl,
            recvPipeOutVec[qpIndex],
            workReqPipeOutVec[qpIndex],
            dmaReadSrvVec[qpIndex],
            dmaWriteSrvVec[qpIndex],
            permCheck4RQ,
            permCheck4SQ,
            pktMetaDataAndPayloadPipeOutVec[idx].reqPktPipeOut,
            pktMetaDataAndPayloadPipeOutVec[idx].respPktPipeOut
        );
        qpDataStreamPipeOutVec[idx] = qp.rdmaReqRespPipeOut;

        // TODO: support CNP
        let addNoErrWorkCompOutRule <- addRules(genEmptyPipeOutRule(
            pktMetaDataAndPayloadPipeOutVec[idx].cnpPipeOut,
            "pktMetaDataAndPayloadPipeOutVec[" + integerToString(idx) +
            "].cnpPipeOut empty assertion @ mkTransportLayerRDMA"
        ));
        // TODO: support CQ
        qpRecvWorkCompPipeOutVec[idx] = qp.workCompPipeOutRQ;
        qpSendWorkCompPipeOutVec[idx] = qp.workCompPipeOutSQ;
    end

    function Bool isDataStreamFinished(DataStream ds) = ds.isLast;
    // TODO: connect to UDP
    let dataStreamPipeOut <- mkPipeOutArbiter(qpDataStreamPipeOutVec, isDataStreamFinished);

    function Bool isWorkCompFinished(WorkComp wc) = True;
    let recvWorkCompPipeOut <- mkPipeOutArbiter(qpRecvWorkCompPipeOutVec, isWorkCompFinished);
    let sendWorkCompPipeOut <- mkPipeOutArbiter(qpSendWorkCompPipeOutVec, isWorkCompFinished);
    let workCompPipeOut <- mkFixedBinaryPipeOutArbiter(
        recvWorkCompPipeOut, sendWorkCompPipeOut
    );

    interface rdmaDataStreamInput   = toPut(inputDataStreamQ);
    interface rdmaDataStreamPipeOut = dataStreamPipeOut;
    interface srvWorkReqRecvReqWorkComp = toGPServer(inputWorkReqOrRecvReqQ, workCompPipeOut);
    interface srvMetaData = metaDataSrv;
endmodule

typedef enum {
    META_DATA_ALLOC_PD,
    META_DATA_CREATE_QP,
    META_DATA_INIT_QP,
    META_DATA_SET_QP_RTR,
    META_DATA_SET_QP_RTS,
    META_DATA_NO_OP
} InitMetaDataState deriving(Bits, Eq, FShow);

module mkInitMetaData#(
    MetaDataSrv metaDataSrv, QpInitAttr qpInitAttr, PipeOut#(AttrQP) qpAttrPipeIn
)(Empty);
    let pdNum = valueOf(MAX_PD);
    let qpNum = valueOf(MAX_QP);
    let qpPerPD = valueOf(TDiv#(MAX_QP, MAX_PD));

    FIFOF#(HandlerPD) pdHandlerQ4Fill <- mkSizedFIFOF(pdNum);
    FIFOF#(QPN)             qpnQ4Init <- mkSizedFIFOF(qpNum);
    FIFOF#(QPN)           qpnQ4Modify <- mkSizedFIFOF(qpNum);

    Count#(Bit#(TLog#(MAX_PD)))                  pdKeyCnt <- mkCount(fromInteger(pdNum - 1));
    Count#(Bit#(TLog#(TAdd#(1, MAX_PD))))        pdReqCnt <- mkCount(fromInteger(pdNum));
    Count#(Bit#(TLog#(MAX_PD)))                 pdRespCnt <- mkCount(fromInteger(pdNum - 1));
    Count#(Bit#(TLog#(TAdd#(1, MAX_QP))))        qpReqCnt <- mkCount(fromInteger(qpNum));
    Count#(Bit#(TLog#(MAX_QP)))                 qpRespCnt <- mkCount(fromInteger(qpNum - 1));
    Count#(Bit#(TLog#(TDiv#(MAX_QP, MAX_PD)))) qpPerPdCnt <- mkCount(fromInteger(qpPerPD - 1));

    Reg#(InitMetaDataState) initMetaDataStateReg <- mkReg(META_DATA_ALLOC_PD);
    // Reg#(Bool)   pdInitDoneReg <- mkReg(False);
    // Reg#(Bool) qpCreateDoneReg <- mkReg(False);
    // Reg#(Bool)   qpInitDoneReg <- mkReg(False);
    // Reg#(Bool) qpModifyDoneReg <- mkReg(False);

    Vector#(MAX_QP, Reg#(Bool)) qpModifyDoneRegVec <- replicateM(mkReg(False));

    // rule reqAllocPDs if (!isZero(pdReqCnt) && !pdInitDoneReg);
    rule reqAllocPDs if (
        !isZero(pdReqCnt) && initMetaDataStateReg == META_DATA_ALLOC_PD
    );
        pdReqCnt.decr(1);

        KeyPD pdKey = zeroExtend(pdKeyCnt);
        pdKeyCnt.incr(1);

        let allocReqPD = ReqPD {
            allocOrNot: True,
            pdKey     : pdKey,
            pdHandler : dontCareValue
        };
        metaDataSrv.request.put(tagged Req4PD allocReqPD);
    endrule

    // rule respAllocPDs if (!pdInitDoneReg);
    rule respAllocPDs if (initMetaDataStateReg == META_DATA_ALLOC_PD);
        if (isZero(pdRespCnt)) begin
            // pdInitDoneReg <= True;
            initMetaDataStateReg <= META_DATA_CREATE_QP;
        end
        else begin
            pdRespCnt.decr(1);
        end

        let maybeAllocRespPD <- metaDataSrv.response.get;
        if (maybeAllocRespPD matches tagged Resp4PD .allocRespPD) begin
            immAssert(
                allocRespPD.successOrNot,
                "allocRespPD.successOrNot assertion @ mkInitMetaData",
                $format(
                    "allocRespPD.successOrNot=", fshow(allocRespPD.successOrNot),
                    " should be true when pdRespCnt=%0d", pdRespCnt
                )
            );
            pdHandlerQ4Fill.enq(allocRespPD.pdHandler);
        end
        else begin
            immFail(
                "maybeAllocRespPD assertion @ mkInitMetaData",
                $format(
                    "maybeAllocRespPD=", fshow(maybeAllocRespPD),
                    " should be Resp4PD"
                )
            );
        end
    endrule

    // rule reqCreateQPs if (!isZero(qpReqCnt) && pdInitDoneReg && !qpCreateDoneReg);
    rule reqCreateQPs if (
        !isZero(qpReqCnt) && initMetaDataStateReg == META_DATA_CREATE_QP
    );
        qpReqCnt.decr(1);

        if (isZero(qpPerPdCnt)) begin
            qpPerPdCnt <= fromInteger(qpPerPD - 1);
            pdHandlerQ4Fill.deq;
        end
        else begin
            qpPerPdCnt.decr(1);
        end

        let pdHandler = pdHandlerQ4Fill.first;

        let createReqQP = ReqQP {
            qpReqType   : REQ_QP_CREATE,
            pdHandler   : pdHandler,
            qpn         : dontCareValue,
            qpAttrMask  : dontCareValue,
            qpAttr      : dontCareValue,
            qpInitAttr  : qpInitAttr
        };
        metaDataSrv.request.put(tagged Req4QP createReqQP);
    endrule

    // rule respCreateQPs if (pdInitDoneReg && !qpCreateDoneReg);
    rule respCreateQPs if (initMetaDataStateReg == META_DATA_CREATE_QP);
        if (isZero(qpRespCnt)) begin
            qpReqCnt  <= fromInteger(qpNum);
            qpRespCnt <= fromInteger(qpNum - 1);
            // qpCreateDoneReg <= True;
            initMetaDataStateReg <= META_DATA_INIT_QP;
        end
        else begin
            qpRespCnt.decr(1);
        end

        let maybeCreateRespQP <- metaDataSrv.response.get;
        if (maybeCreateRespQP matches tagged Resp4QP .createRespQP) begin
            immAssert(
                createRespQP.successOrNot,
                "createRespQP.successOrNot assertion @ mkInitMetaData",
                $format(
                    "createRespQP.successOrNot=", fshow(createRespQP.successOrNot),
                    " should be true when qpRespCnt=%0d", qpRespCnt
                )
            );

            let qpn = createRespQP.qpn;
            qpnQ4Init.enq(qpn);
            // $display(
            //     "time=%0t: createRespQP=", $time, fshow(createRespQP),
            //     " should be success, and qpn=%h, qpRespCnt=%h",
            //     qpn, qpRespCnt
            // );
        end
        else begin
            immFail(
                "maybeCreateRespQP assertion @ mkInitMetaData",
                $format(
                    "maybeCreateRespQP=", fshow(maybeCreateRespQP),
                    " should be Resp4QP"
                )
            );
        end
    endrule

    // rule reqInitQPs if (
    //     !isZero(qpReqCnt) &&
    //     pdInitDoneReg     &&
    //     qpCreateDoneReg   &&
    //     !qpInitDoneReg
    // );
    rule reqInitQPs if (
        !isZero(qpReqCnt) && initMetaDataStateReg == META_DATA_INIT_QP
    );
        qpReqCnt.decr(1);

        let qpn = qpnQ4Init.first;
        qpnQ4Init.deq;

        let qpAttr = qpAttrPipeIn.first;
        qpAttr.qpState = IBV_QPS_INIT;
        let initReqQP = ReqQP {
            qpReqType   : REQ_QP_MODIFY,
            pdHandler   : dontCareValue,
            qpn         : qpn,
            qpAttrMask  : getReset2InitRequiredAttr,
            qpAttr      : qpAttr,
            qpInitAttr  : dontCareValue
        };
        metaDataSrv.request.put(tagged Req4QP initReqQP);
    endrule

    // rule respInitQPs if (pdInitDoneReg && qpCreateDoneReg && !qpInitDoneReg);
    rule respInitQPs if (initMetaDataStateReg == META_DATA_INIT_QP);
        if (isZero(qpRespCnt)) begin
            qpReqCnt  <= fromInteger(qpNum);
            qpRespCnt <= fromInteger(qpNum - 1);
            // qpInitDoneReg <= True;
            initMetaDataStateReg <= META_DATA_SET_QP_RTR;
        end
        else begin
            qpRespCnt.decr(1);
        end

        let maybeInitRespQP <- metaDataSrv.response.get;
        if (maybeInitRespQP matches tagged Resp4QP .initRespQP) begin
            immAssert(
                initRespQP.successOrNot,
                "initRespQP.successOrNot assertion @ mkInitMetaData",
                $format(
                    "initRespQP.successOrNot=", fshow(initRespQP.successOrNot),
                    " should be true when qpRespCnt=%0d", qpRespCnt
                )
            );

            let qpn = initRespQP.qpn;
            qpnQ4Modify.enq(qpn);
            // $display(
            //     "time=%0t: initRespQP=", $time, fshow(initRespQP),
            //     " should be success, and qpn=%h, qpRespCnt=%h",
            //     $time, qpn, qpRespCnt
            // );
        end
        else begin
            immFail(
                "maybeInitRespQP assertion @ mkInitMetaData",
                $format(
                    "maybeInitRespQP=", fshow(maybeInitRespQP),
                    " should be Resp4QP"
                )
            );
        end
    endrule

    // rule reqModifyQPs if (
    //     !isZero(qpReqCnt) &&
    //     pdInitDoneReg     &&
    //     qpCreateDoneReg   &&
    //     qpInitDoneReg     &&
    //     !qpModifyDoneReg
    // );
    rule reqRtrQPs if (
        !isZero(qpReqCnt) && initMetaDataStateReg == META_DATA_SET_QP_RTR
    );
        qpReqCnt.decr(1);

        let qpn = qpnQ4Modify.first;
        qpnQ4Modify.deq;

        let qpAttr = qpAttrPipeIn.first;
        qpAttrPipeIn.deq;

        qpAttr.qpState = IBV_QPS_RTR;
        let setRtrReqQP = ReqQP {
            qpReqType   : REQ_QP_MODIFY,
            pdHandler   : dontCareValue,
            qpn         : qpn,
            qpAttrMask  : getInit2RtrRequiredAttr,
            qpAttr      : qpAttr,
            qpInitAttr  : dontCareValue
        };
        metaDataSrv.request.put(tagged Req4QP setRtrReqQP);
    endrule

    // rule respModifyQPs if (
    //     pdInitDoneReg   &&
    //     qpCreateDoneReg &&
    //     qpInitDoneReg   &&
    //     !qpModifyDoneReg
    // );
    rule respRtrQPs if (initMetaDataStateReg == META_DATA_SET_QP_RTR);
        if (isZero(qpRespCnt)) begin
            // qpModifyDoneReg <= True;
            initMetaDataStateReg <= META_DATA_SET_QP_RTS;
        end
        else begin
            qpRespCnt.decr(1);
        end

        let maybeModifyRespQP <- metaDataSrv.response.get;
        if (maybeModifyRespQP matches tagged Resp4QP .setRtrRespQP) begin
            immAssert(
                setRtrRespQP.successOrNot,
                "setRtrRespQP.successOrNot assertion @ mkInitMetaData",
                $format(
                    "setRtrRespQP.successOrNot=", fshow(setRtrRespQP.successOrNot),
                    " should be true when qpRespCnt=%0d", qpRespCnt,
                    ", setRtrRespQP=", fshow(setRtrRespQP)
                )
            );
            // $display(
            //     "time=%0t: setRtrRespQP=", $time, fshow(setRtrRespQP),
            //     " should be success, and setRtrRespQP.qpn=%h, qpRespCnt=%h",
            //     $time, setRtrRespQP.qpn, qpRespCnt
            // );
        end
        else begin
            immFail(
                "maybeModifyRespQP assertion @ mkInitMetaData",
                $format(
                    "maybeModifyRespQP=", fshow(maybeModifyRespQP),
                    " should be Resp4QP"
                )
            );
        end
    endrule

    // rule reqModifyQPs if (
    //     !isZero(qpReqCnt) &&
    //     pdInitDoneReg     &&
    //     qpCreateDoneReg   &&
    //     qpInitDoneReg     &&
    //     !qpModifyDoneReg
    // );
    rule reqRtsQPs if (
        !isZero(qpReqCnt) && initMetaDataStateReg == META_DATA_SET_QP_RTS
    );
        qpReqCnt.decr(1);

        let qpn = qpnQ4Modify.first;
        qpnQ4Modify.deq;

        let qpAttr = qpAttrPipeIn.first;
        qpAttrPipeIn.deq;

        qpAttr.qpState = IBV_QPS_RTS;
        let setRtsReqQP = ReqQP {
            qpReqType   : REQ_QP_MODIFY,
            pdHandler   : dontCareValue,
            qpn         : qpn,
            qpAttrMask  : getRtr2RtsRequiredAttr,
            qpAttr      : qpAttr,
            qpInitAttr  : dontCareValue
        };
        metaDataSrv.request.put(tagged Req4QP setRtsReqQP);
    endrule

    // rule respModifyQPs if (
    //     pdInitDoneReg   &&
    //     qpCreateDoneReg &&
    //     qpInitDoneReg   &&
    //     !qpModifyDoneReg
    // );
    rule respRtsQPs if (initMetaDataStateReg == META_DATA_SET_QP_RTS);
        if (isZero(qpRespCnt)) begin
            // qpModifyDoneReg <= True;
            initMetaDataStateReg <= META_DATA_NO_OP;
        end
        else begin
            qpRespCnt.decr(1);
        end

        let maybeModifyRespQP <- metaDataSrv.response.get;
        if (maybeModifyRespQP matches tagged Resp4QP .setRtsRespQP) begin
            immAssert(
                setRtsRespQP.successOrNot,
                "setRtsRespQP.successOrNot assertion @ mkInitMetaData",
                $format(
                    "setRtsRespQP.successOrNot=", fshow(setRtsRespQP.successOrNot),
                    " should be true when qpRespCnt=%0d", qpRespCnt,
                    ", setRtsRespQP=", fshow(setRtsRespQP)
                )
            );
            // $display(
            //     "time=%0t: setRtsRespQP=", $time, fshow(setRtsRespQP),
            //     " should be success, and setRtsRespQP.qpn=%h, qpRespCnt=%h",
            //     $time, setRtsRespQP.qpn, qpRespCnt
            // );
        end
        else begin
            immFail(
                "maybeModifyRespQP assertion @ mkInitMetaData",
                $format(
                    "maybeModifyRespQP=", fshow(maybeModifyRespQP),
                    " should be Resp4QP"
                )
            );
        end
    endrule
endmodule

// TODO: connect to DMA IP

// This function should be used in simulation only
function Tuple3#(TotalFragNum, ByteEn, ByteEnBitNum) calcTotalFragNumByLength(Length dmaLen);
    Bit#(DATA_BUS_BYTE_NUM_WIDTH) lastFragByteNumResidue = truncate(dmaLen);
    Bit#(TSub#(RDMA_MAX_LEN_WIDTH, DATA_BUS_BYTE_NUM_WIDTH)) truncatedLen = truncateLSB(dmaLen);
    let lastFragEmpty = isZero(lastFragByteNumResidue);
    TotalFragNum fragNum = zeroExtend(truncatedLen + zeroExtend(pack(!lastFragEmpty)));

    // let shiftAmt = valueOf(TLog#(DATA_BUS_BYTE_WIDTH));
    // TotalFragNum fragNum = truncate(dmaLen >> shiftAmt);
    // BusByteWidthMask busByteWidthMask = maxBound;
    // let lastFragSize = truncate(dmaLen) & busByteWidthMask;
    // Bool lastFragEmpty = isZero(lastFragSize);
    // if (!lastFragEmpty) begin
    //     fragNum = fragNum + 1;
    // end

    ByteEnBitNum lastFragValidByteNum = lastFragEmpty ?
        fromInteger(valueOf(DATA_BUS_BYTE_WIDTH)) :
        zeroExtend(lastFragByteNumResidue);
    ByteEn lastFragByteEn = genByteEn(lastFragValidByteNum);
    return tuple3(fragNum, lastFragByteEn, lastFragValidByteNum);
endfunction

module mkDmaReadSrv(DmaReadSrv);
    FIFOF#(DmaReadReq) dmaReadReqQ <- mkFIFOF;
    FIFOF#(DmaReadResp) dmaReadRespQ <- mkFIFOF;

    Reg#(TotalFragNum) totalFragCntReg <- mkRegU;
    Reg#(Bool) busyReg <- mkReg(False);
    Reg#(Bool) isFirstReg <- mkRegU;
    Reg#(ByteEn) lastFragByteEnReg <- mkRegU;
    Reg#(BusBitNum) lastFragInvalidBitNumReg <- mkRegU;
    Reg#(DmaReadReq) curReqReg <- mkRegU;

    Bool isFragCntZero = isZero(totalFragCntReg);

    rule acceptReq if (!busyReg);
        let curReq = dmaReadReqQ.first;
        dmaReadReqQ.deq;

        let isZeroLen = isZero(curReq.len);
        immAssert(
            !isZeroLen,
            "dmaReadReq.len non-zero assrtion",
            $format("curReq.len=%h should not be zero", curReq.len)
        );

        let { totalFragCnt, lastFragByteEn, lastFragValidByteNum } =
            calcTotalFragNumByLength(curReq.len);
        let { lastFragValidBitNum, lastFragInvalidByteNum, lastFragInvalidBitNum } =
            calcFragBitNumAndByteNum(lastFragValidByteNum);

        totalFragCntReg <= isZeroLen ? 0 : totalFragCnt - 1;
        lastFragByteEnReg <= lastFragByteEn;
        lastFragInvalidBitNumReg <= lastFragInvalidBitNum;

        immAssert(
            !isZero(lastFragByteEn),
            "lastFragByteEn non-zero assertion",
            $format(
                "lastFragByteEn=%h should not have zero ByteEn, curReq.len=%h",
                lastFragByteEn, curReq.len
            )
        );

        curReqReg <= curReq;
        busyReg <= True;
        isFirstReg <= True;

        // $display(
        //     "time=%0t: curReq.len=%0d, totalFragCnt=%0d",
        //     $time, curReq.len, totalFragCnt
        // );
    endrule

    rule genResp if (busyReg);
        totalFragCntReg <= totalFragCntReg - 1;
        DataStream dataStream = dontCareValue;
        dataStream.isFirst = isFirstReg;
        isFirstReg <= False;
        dataStream.isLast = isFragCntZero;
        dataStream.byteEn = maxBound;

        if (isFragCntZero) begin
            busyReg <= False;
            dataStream.byteEn = lastFragByteEnReg;
            DATA tmpData = dataStream.data >> lastFragInvalidBitNumReg;
            dataStream.data = truncate(tmpData << lastFragInvalidBitNumReg);
        end

        let resp = DmaReadResp {
            initiator : curReqReg.initiator,
            sqpn      : curReqReg.sqpn,
            wrID      : curReqReg.wrID,
            isRespErr : False,
            dataStream: dataStream
        };
        dmaReadRespQ.enq(resp);

        immAssert(
            !isZero(dataStream.byteEn),
            "dmaReadResp.data.byteEn non-zero assertion",
            $format("dmaReadResp.data should not have zero ByteEn, ", fshow(dataStream))
        );
        // $display(
        //     "time=%0t: mkSimDmaReadSrvAndReqRespPipeOut response, totalFragNum=%h, dataStream=",
        //     $time, totalFragCntReg, fshow(dataStream)
        // );
    endrule

    return toGPServer(dmaReadReqQ, dmaReadRespQ);
endmodule

module mkDmaWriteSrv(DmaWriteSrv);
    FIFOF#(DmaWriteReq) dmaWriteReqQ <- mkFIFOF;
    FIFOF#(DmaWriteResp) dmaWriteRespQ <- mkFIFOF;

    function Action genDmaWriteResp(DmaWriteMetaData metaData);
        action
            let dmaWriteResp = DmaWriteResp {
                initiator: metaData.initiator,
                sqpn     : metaData.sqpn,
                psn      : metaData.psn,
                isRespErr: False
            };
            // $display("time=%0t: dmaWriteResp=", $time, fshow(dmaWriteResp));

            dmaWriteRespQ.enq(dmaWriteResp);
        endaction
    endfunction

    rule write;
        let dmaWriteReq = dmaWriteReqQ.first;
        dmaWriteReqQ.deq;

        // $display("time=%0t: dmaWriteReq=", $time, fshow(dmaWriteReq));

        if (dmaWriteReq.dataStream.isLast) begin
            genDmaWriteResp(dmaWriteReq.metaData);
        end
    endrule

    return toGPServer(dmaWriteReqQ, dmaWriteRespQ);
endmodule
