// Adjustible settings
typedef 32 MAX_PENDING_REQ_NUM;
// typedef 16 MAX_PENDING_READ_ATOMIC_REQ_NUM;
typedef 256 DATA_BUS_WIDTH;
typedef TExp#(31) MAX_MR_SIZE; // 2GB
